package environment_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import item_pack::*;
  import sequence_pack::*;

  import input_agent_pack::*;
  import output_agent_pack::*;

  `include "src/test/environment/coverage/input_covergroup.sv"
  `include "src/test/environment/coverage/output_covergroup.sv" 

  `include "src/test/environment/coverage/coverage.svh"

  `include "src/test/environment/virtual_sequencer.svh"
  `include "src/test/sequence/virtual_sequence.svh"
  
  `include "src/test/environment/environment_config.svh"
  `include "src/test/environment/environment.svh"
endpackage : environment_pack