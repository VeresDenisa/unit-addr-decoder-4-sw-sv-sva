package environment_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import item_pack::*;
  import sequence_pack::*;

  import input_agent_pack::*;
  import output_agent_pack::*;

  import coverage_pack::*;

  `include "src/test/environment/virtual_sequencer.svh"
  `include "src/test/environment/environment_config.svh"
  `include "src/test/environment/environment.svh"
endpackage : environment_pack