package input_agent_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  import item_pack::*;

  `include "src/test/environment/input_agent/input_config.svh"

  `include "src/test/environment/input_agent/input_driver.svh"
  `include "src/test/environment/input_agent/input_monitor.svh"
  
  `include "src/test/environment/input_agent/input_agent.svh"
endpackage : input_agent_pack