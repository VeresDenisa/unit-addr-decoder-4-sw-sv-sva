package test_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import item_pack::*;
  import sequence_pack::*;

  import environment_pack::*;

  `include "src/test/test.svh"
endpackage : test_pack