package sequence_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import item_pack::*;

  `include "src/test/sequence/input_sequence.svh"
  `include "src/test/sequence/output_sequence.svh"
endpackage : sequence_pack