package coverage_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "src/test/environment/coverage/input_covergroup.sv"
  `include "src/test/environment/coverage/output_covergroup.sv" 

  `include "src/test/environment/coverage/coverage.svh"
endpackage : coverage_pack