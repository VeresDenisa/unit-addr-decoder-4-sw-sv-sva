package item_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "src/test/item/input_item.svh"
  `include "src/test/item/output_item.svh"
endpackage : item_pack