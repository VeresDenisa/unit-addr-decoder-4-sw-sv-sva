package output_agent_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "src/test/environment/output_agent/output_config.svh"

  `include "src/test/environment/output_agent/output_sequencer.svh"
  `include "src/test/environment/output_agent/output_driver.svh"
  `include "src/test/environment/output_agent/output_monitor.svh"
  
  `include "src/test/environment/output_agent/output_agent.svh"
endpackage : output_agent_pack